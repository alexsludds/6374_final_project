/afs/athena.mit.edu/dept/cadence/GPDK045/gsclib045_all_v4.4/gsclib045/lef/gsclib045_tech.lef